`define RESET 3'b001
`define IDLE  3'b010
`define START 3'b011
`define DATA  3'b100
`define PARITY 3'b101
`define STOP  3'b110
